module Shifter (
    leftRight,
    shamt,
    sftSrc,
    result
);

  //I/O ports
  input leftRight;        //1 bit
  input [5-1:0] shamt;    //5 bits
  input [32-1:0] sftSrc;  //32 bits

  output [32-1:0] result; //32 bits

  //Internal Signals
  wire [32-1:0] result;



  //Main function
  /*your code here*/
assign result = (~leftRight) ? (sftSrc << shamt) : (sftSrc >> shamt);


endmodule
